`ifndef _io_params_vh_
`define _io_params_vh_
parameter _CLK_PER_HALF_BIT = 20;
`endif