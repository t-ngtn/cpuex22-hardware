`ifndef _params_vh_
`define _params_vh_

`endif