// 各値の定義
// 使わなかった、、