// 各値の定義

// Core全体

// ALU

// ControlUnit

// RegFile

// InstMem

// 